
package comp1_env1_test_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    
    import comp1_env1_env_pkg::*;

    `include "comp1_test_utils.svh"
    `include "env1_base_test.svh"

endpackage