
module comp1_env1_wrapper (comp1_env1_tb_if tb_if);

    // connect DUT here

endmodule
