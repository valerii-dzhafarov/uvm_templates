package comp1_env1_env_pkg;

    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "env1_cfg.svh"
    `include "env1_env.svh"

endpackage