package comp1_env1_env_pkg;

    import uvm_pkg::*;
    `include "uvm_macros.svh"


    import comp1_agent1_pkg::*; // ut_del_pragma
    `include "stack_model.svh"  // ut_del_pragma
    `include "env1_stack_sb.svh"  // ut_del_pragma

    `include "env1_cfg.svh"
    `include "env1_env.svh"
endpackage