
module inst_test;

    import comp1_agent1_pkg::*;
    comp1_agent1_if agent1_if(1,1);

endmodule