interface comp1_env1_tb_if;

endinterface
