package comp1_agent1_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "agent1_config.svh"
    `include "agent1_item.svh"

    `include "agent1_driver.svh"
    `include "agent1_monitor.svh"
    `include "agent1_sequencer.svh"

    `include "agent1_checker.svh"
    `include "agent1_cov_collector.svh"

    `include "agent1_agent.svh"

    `include "agent1_base_seq.svh"
endpackage